module sync_apb2core (
    
);


endmodule