module apb_slave_interface (
    ports
);
    
endmodule