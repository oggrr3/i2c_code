`ifdef SCOREBOARD 
`define SCOREBOARD

    class scoreboard;
        bit         sda         ;
        bit [7:0]   prdata      ;

    endclass

`endif macro